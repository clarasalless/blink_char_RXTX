`timescale 1ns/1ps
module
CoreTimer
(
PCLK
,
PRESETn
,
PENABLE
,
PSEL
,
PADDR
,
PWRITE
,
PWDATA
,
PRDATA
,
TIMINT
)
;
`define CoreTimer_O  \
3 \
'b \
000
`define CoreTimer_I  \
3 \
'b \
001
`define CoreTimer_l  \
3 \
'b \
010
`define CoreTimer_OI  \
3 \
'b \
011
`define CoreTimer_II  \
3 \
'b \
100
`define CoreTimer_lI  \
3 \
'b \
101
`define CoreTimer_Ol  \
3 \
'b \
110
parameter
WIDTH
=
32
;
parameter
INTACTIVEH
=
1
;
input
PCLK
;
input
PRESETn
;
input
PENABLE
;
input
PSEL
;
input
[
4
:
2
]
PADDR
;
input
PWRITE
;
input
[
31
:
0
]
PWDATA
;
output
[
31
:
0
]
PRDATA
;
output
TIMINT
;
wire
PCLK
;
wire
PRESETn
;
wire
PENABLE
;
wire
[
4
:
2
]
PADDR
;
wire
PWRITE
;
wire
[
31
:
0
]
PWDATA
;
wire
[
31
:
0
]
PRDATA
;
wire
PSEL
;
wire
TIMINT
;
wire
[
31
:
0
]
CoreTimer_Il
;
reg
[
31
:
0
]
CoreTimer_ll
;
wire
CoreTimer_O0
;
reg
[
31
:
0
]
CoreTimer_I0
;
wire
CoreTimer_l0
;
reg
[
6
:
0
]
CoreTimer_O1
;
wire
CoreTimer_I1
;
wire
CoreTimer_l1
;
wire
CoreTimer_OOI
;
wire
CoreTimer_IOI
;
wire
CoreTimer_lOI
;
wire
CoreTimer_OII
;
reg
[
3
:
0
]
CoreTimer_III
;
wire
CoreTimer_lII
;
reg
CoreTimer_OlI
;
reg
[
WIDTH
-
1
:
0
]
CoreTimer_IlI
;
reg
[
9
:
0
]
CoreTimer_llI
;
reg
[
WIDTH
-
1
:
0
]
CoreTimer_O0I
;
wire
CoreTimer_I0I
;
reg
CoreTimer_l0I
;
wire
CoreTimer_O1I
;
reg
CoreTimer_I1I
;
wire
CoreTimer_l1I
;
wire
CoreTimer_OOl
;
reg
CoreTimer_IOl
;
wire
CoreTimer_lOl
;
reg
CoreTimer_OIl
;
reg
CoreTimer_IIl
;
assign
CoreTimer_l0
=
(
PADDR
==
`CoreTimer_l
)
?
(
PWRITE
&&
PSEL
&&
!
PENABLE
)
:
1
'b
0
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_lIl
if
(
!
PRESETn
)
CoreTimer_O1
<=
3
'b
000
;
else
if
(
CoreTimer_l0
)
CoreTimer_O1
<=
PWDATA
[
2
:
0
]
;
end
assign
CoreTimer_I1
=
CoreTimer_O1
[
2
]
;
assign
CoreTimer_l1
=
CoreTimer_O1
[
1
]
;
assign
CoreTimer_OOI
=
CoreTimer_O1
[
0
]
;
assign
CoreTimer_IOI
=
(
CoreTimer_I1
==
1
'b
1
)
?
1
'b
1
:
1
'b
0
;
assign
CoreTimer_lOI
=
CoreTimer_OOl
&&
CoreTimer_IOI
&&
(
CoreTimer_l0
&&
!
PWDATA
[
2
]
)
;
assign
CoreTimer_OII
=
(
PADDR
==
`CoreTimer_OI
)
?
(
PWRITE
&&
PSEL
&&
!
PENABLE
)
:
1
'b
0
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_Oll
if
(
!
PRESETn
)
CoreTimer_III
<=
4
'b
0000
;
else
if
(
CoreTimer_OII
)
CoreTimer_III
<=
PWDATA
[
3
:
0
]
;
end
assign
CoreTimer_lII
=
(
PADDR
==
`CoreTimer_O
)
?
(
PWRITE
&&
PSEL
&&
!
PENABLE
)
:
1
'b
0
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_Ill
if
(
!
PRESETn
)
CoreTimer_OlI
<=
1
'b
0
;
else
CoreTimer_OlI
<=
CoreTimer_lII
;
end
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_lll
if
(
!
PRESETn
)
CoreTimer_IlI
<=
{
WIDTH
{
1
'b
0
}
}
;
else
if
(
CoreTimer_lII
)
CoreTimer_IlI
<=
PWDATA
[
WIDTH
-
1
:
0
]
;
end
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_O0l
if
(
!
PRESETn
)
CoreTimer_llI
<=
{
10
{
1
'b
0
}
}
;
else
if
(
CoreTimer_OlI
||
CoreTimer_lOI
)
CoreTimer_llI
<=
{
10
{
1
'b
0
}
}
;
else
CoreTimer_llI
<=
CoreTimer_llI
+
1
'b
1
;
end
always
@
(
CoreTimer_llI
or
CoreTimer_III
)
begin
:
CoreTimer_I0l
CoreTimer_IIl
=
1
'b
0
;
case
(
CoreTimer_III
)
4
'b
0000
:
if
(
CoreTimer_llI
[
0
]
==
1
'b
1
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
0001
:
if
(
CoreTimer_llI
[
1
:
0
]
==
2
'b
11
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
0010
:
if
(
CoreTimer_llI
[
2
:
0
]
==
3
'b
111
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
0011
:
if
(
CoreTimer_llI
[
3
:
0
]
==
4
'b
1111
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
0100
:
if
(
CoreTimer_llI
[
4
:
0
]
==
5
'b
11111
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
0101
:
if
(
CoreTimer_llI
[
5
:
0
]
==
6
'b
111111
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
0110
:
if
(
CoreTimer_llI
[
6
:
0
]
==
7
'b
1111111
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
0111
:
if
(
CoreTimer_llI
[
7
:
0
]
==
8
'b
11111111
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
1000
:
if
(
CoreTimer_llI
[
8
:
0
]
==
9
'b
111111111
)
CoreTimer_IIl
=
1
'b
1
;
4
'b
1001
:
if
(
CoreTimer_llI
[
9
:
0
]
==
10
'b
1111111111
)
CoreTimer_IIl
=
1
'b
1
;
default
:
if
(
CoreTimer_llI
[
9
:
0
]
==
10
'b
1111111111
)
CoreTimer_IIl
=
1
'b
1
;
endcase
end
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_l0l
if
(
!
PRESETn
)
CoreTimer_OIl
<=
1
'b
0
;
else
CoreTimer_OIl
<=
CoreTimer_IIl
;
end
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_O1l
if
(
!
PRESETn
)
CoreTimer_O0I
<=
{
WIDTH
{
1
'b
1
}
}
;
else
if
(
CoreTimer_OlI
||
CoreTimer_lOI
)
CoreTimer_O0I
<=
CoreTimer_IlI
;
else
if
(
CoreTimer_OOI
&&
CoreTimer_OIl
)
if
(
CoreTimer_OOl
)
if
(
CoreTimer_IOI
)
CoreTimer_O0I
<=
CoreTimer_O0I
;
else
CoreTimer_O0I
<=
CoreTimer_IlI
;
else
CoreTimer_O0I
<=
CoreTimer_O0I
-
1
'b
1
;
end
assign
CoreTimer_OOl
=
(
CoreTimer_O0I
==
{
WIDTH
{
1
'b
0
}
}
)
?
1
'b
1
:
1
'b
0
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_I1l
if
(
!
PRESETn
)
CoreTimer_IOl
<=
1
'b
0
;
else
CoreTimer_IOl
<=
CoreTimer_OOl
;
end
assign
CoreTimer_lOl
=
CoreTimer_OOl
&&
!
CoreTimer_IOl
;
assign
CoreTimer_O1I
=
(
CoreTimer_lOl
||
CoreTimer_I1I
)
&&
(
!
CoreTimer_l0I
)
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_l1l
if
(
!
PRESETn
)
CoreTimer_I1I
<=
1
'b
0
;
else
CoreTimer_I1I
<=
CoreTimer_O1I
;
end
assign
CoreTimer_l1I
=
CoreTimer_I1I
&&
CoreTimer_l1
;
assign
TIMINT
=
(
INTACTIVEH
)
?
CoreTimer_l1I
:
!
CoreTimer_l1I
;
assign
CoreTimer_I0I
=
(
PADDR
==
`CoreTimer_II
)
?
(
PWRITE
&&
PSEL
&&
!
PENABLE
)
:
1
'b
0
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_OO0
if
(
!
PRESETn
)
CoreTimer_l0I
<=
1
'b
0
;
else
if
(
CoreTimer_I0I
)
CoreTimer_l0I
<=
1
'b
1
;
else
CoreTimer_l0I
<=
1
'b
0
;
end
always
@
(
PWRITE
or
PSEL
or
PADDR
or
CoreTimer_IlI
or
CoreTimer_O0I
or
CoreTimer_O1
or
CoreTimer_III
or
CoreTimer_I1I
or
CoreTimer_l1I
)
begin
:
CoreTimer_IO0
CoreTimer_I0
=
{
32
{
1
'b
0
}
}
;
if
(
!
PWRITE
&&
PSEL
)
case
(
PADDR
)
`CoreTimer_O
:
CoreTimer_I0
[
WIDTH
-
1
:
0
]
=
CoreTimer_IlI
;
`CoreTimer_I
:
CoreTimer_I0
[
WIDTH
-
1
:
0
]
=
CoreTimer_O0I
;
`CoreTimer_l
:
CoreTimer_I0
[
2
:
0
]
=
CoreTimer_O1
;
`CoreTimer_OI
:
CoreTimer_I0
[
3
:
0
]
=
CoreTimer_III
;
`CoreTimer_lI
:
CoreTimer_I0
[
0
]
=
CoreTimer_I1I
;
`CoreTimer_Ol
:
CoreTimer_I0
[
0
]
=
CoreTimer_l1I
;
default
:
CoreTimer_I0
=
{
32
{
1
'b
0
}
}
;
endcase
else
CoreTimer_I0
=
{
32
{
1
'b
0
}
}
;
end
assign
CoreTimer_O0
=
(
PSEL
&&
!
PWRITE
&&
!
PENABLE
)
;
assign
CoreTimer_Il
=
(
CoreTimer_O0
)
?
CoreTimer_I0
:
{
32
{
1
'b
0
}
}
;
always
@
(
negedge
PRESETn
or
posedge
PCLK
)
begin
:
CoreTimer_lO0
if
(
!
PRESETn
)
CoreTimer_ll
<=
{
32
{
1
'b
0
}
}
;
else
CoreTimer_ll
<=
CoreTimer_Il
;
end
assign
PRDATA
=
CoreTimer_ll
;
endmodule
